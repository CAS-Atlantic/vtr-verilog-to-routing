module simple_op(out,a,b);
input a;
input b;
output out;

xnor(out,a,b);
endmodule 