//And 
module simple_op(a,b,out);
    input a;
    input b;
    output out;

    and(out,a,b);
endmodule

