module simple_op(out,a,b);
input a;
input b;
output out;

nand(out,a,b);
endmodule 
