module simple_op(a,b,out);
input a;
input b;
output out;

or(out,a,b);
endmodule 