module simple_op(out,a,b);
input a;
input b;
output out;

xor(out,a,b);
endmodule 