module simple_op(a, out);
    input   a;
    output  out;

    not(out, a);
endmodule