//And 
module simple_op(a,b,c,d,out);
    input a;
    input b;
    input c;
    input d;
    output out;

    and(out,a,b,c,d);
endmodule

