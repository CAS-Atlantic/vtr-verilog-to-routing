module simple_op(out,a,b);
input a;
input b;
output out;

nor(out,a,b);
endmodule 